  module backtrack_unit(input logic backtrack,
                      input logic ,)
					  
					  
					  
  endmodule					  