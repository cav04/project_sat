module main;
initial $hello;
initial #100 $linkc;
initial #200 $linkc;
endmodule