module mux_8_1(
			input logic input1,
				input logic input1,)